module dot(ctrl,key,clk,led_r,led_g,row);
input [2:0]ctrl;
input [6:0]key;
input clk;
output reg [7:0]led_r;
output reg [7:0]led_g;
output reg [7:0]row;

parameter d=2000;
reg i=4'd4999;
reg [2:0]cnt=3'b000;
always @(posedge clk) begin
if(cnt==3'b111)
	cnt<=3'b000;
else cnt=cnt+1'b1;
end
always @(*)begin
	/*if(ctrl==3'b100)begin*/
 case(cnt)
 3'b000:begin led_r[7:0]=8'b0000_0001;
	led_g[7:0]=8'b0000_0001;
	row[7:0]=8'b1111_1110;end

 3'b001:begin led_r[7:0]=8'b0000_0010;
	led_g[7:0]=8'b0000_0010;
	row[7:0]=8'b1111_1100;end
	
 3'b010:begin led_r[7:0]=8'b0000_0100;
	led_g[7:0]=8'b0000_0100;
	row[7:0]=8'b1111_1000;end
	
 3'b011:begin led_r[7:0]=8'b0000_1000;
	led_g[7:0]=8'b0000_1000;
	row[7:0]=8'b1111_0000;end
	
 3'b100:begin led_r[7:0]=8'b0001_0000;
	led_g[7:0]=8'b0001_0000;
	row[7:0]=8'b1110_0000;end
	
 3'b101:begin led_r[7:0]=8'b0010_0000;
	led_g[7:0]=8'b0010_0000;
	row[7:0]=8'b1100_0000;end
	
 3'b110:begin led_r[7:0]=8'b0100_0000;
	led_g[7:0]=8'b0100_0000;
	row[7:0]=8'b1000_0000;end
	
 3'b111:begin led_r[7:0]=8'b0000_0000;
	led_g[7:0]=8'b0000_0000;
	row[7:0]=8'b0000_0000;end
endcase
	//end*/
end

endmodule 

module play();
endmodule 

module auto_play();
endmodule 
